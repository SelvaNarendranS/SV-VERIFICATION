// interface 

interface intf;
  
  logic clk;
  logic reset;
  logic d;
  logic q;
  logic q_bar;
  
endinterface